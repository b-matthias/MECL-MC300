MC306.cir
*
* SPICE netlist for the Motorola MC306 ECL circuit
*
* Expandable 3-input gate, output OR and NOR
* see also MC307 and MC305
* ref page 2-9
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC306 vbb vee vcc or nor in1 in2 in3 ehi elo
*             1   2   3   4  5   6   7   8   9   10
rc1    vcc     ehi             290
rc2    vcc     n02             315
q1     ehi     in1     elo     2N3904
q2     ehi     in2     elo     2N3904
q3     ehi     in3     elo     2N3904
q4     n02     vbb     elo     2N3904
re1    elo     vee             1240
q5     vcc     ehi     nor     2N3904
q6     vcc     n02     or      2N3904
ro1    nor     vee             2000
ro2    or      vee             2000
.ends MC306

.end
