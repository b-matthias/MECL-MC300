MC301.cir
*
* SPICE netlist for the Motorola MC301 ECL circuit
*
*  5-input gate, output OR and NOR
* ref page 2-9
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC301 vbb  vee  vcc  or nor in1 in2 in3 in4 in5
*             vbb  vee  vcc  tp
rc1    vcc     n01             290
rc2    vcc     n02             315
q1     n01     in1     n03     2N3904
q2     n01     in2     n03     2N3904
q3     n01     in3     n03     2N3904
q4     n01     in4     n03     2N3904
q5     n01     in5     n03     2N3904
q6     n02     vbb     n03     2N3904
re1    n03     vee             1240
q7     vcc     n01     nor     2N3904
q8     vcc     n02     or      2N3904
ro1    nor     vee             2000
ro2    or      vee             2000
.ends MC301

.end
