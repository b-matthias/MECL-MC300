MC352A.cir
*
* SPICE netlist for the Motorola MC352A ECL circuit
*
* R-S Flip-Flop, DC coupled with expandable input
* ref page 2-52
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC352A ehi vee vcc nq q set1 set2 elo res1 res2
*             1   2   3   4  5 6    7    8   9    10
rc1    vcc     n01             220
rc2    vcc     ehi             220
q1     vcc     n01     nq      2N3904
q2     vcc     n01     n02     2N3904
q3     vcc     ehi     n03     2N3904
q4     vcc     ehi     q       2N3904
q5     n01     set1    elo     2N3904
q6     n01     set2    elo     2N3904
q7     n01     n03     n04     2N3904
q8     ehi     n02     n04     2N3904
q9     ehi     res1    elo     2N3904
q10    ehi     res2    elo     2N3904
ro1    nq      vee             2000
re1    n02     elo             2400
re2    n04     elo             75
re3    elo     vee             875
re4    n03     elo             2400
ro2    q       vee             2000
.ends MC352A

.end
