MC307.cir
*
* SPICE netlist for the Motorola MC307 ECL circuit
*
* Expandable 3-input gate, output OR and NOR
* see also MC306
* ref page 2-9
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC307 vbb  vee  vcc or nor in1 in2 in3 exphi explo
*             vbb  vee  vcc  tp
rc1    vcc     exphi           290
rc2    vcc     n02             315
q1     exphi   in1     explo   2N3904
q2     exphi   in2     explo   2N3904
q3     exphi   in3     explo   2N3904
q4     n02     vbb     explo   2N3904
re1    explo   vee             1240
q5     vcc     exphi   nor     2N3904
q6     vcc     n02     or      2N3904
.ends MC307

.end
