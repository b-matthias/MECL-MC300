MC312A.cir
*
* SPICE netlist for the Motorola MC312A ECL circuit
*
* Dual 2-input gates, output NOR
* see also MC312G.cir, MC312F.cir and MC312.md
* ref page 2-16
*
* Models
*
.import 2N3904.mod
.import 1N4148.mod
*
* Circuit netlist
*
.subckt MC312A in6 vee vcc nor2 nor1 in1 in2 in3 in4 in5
*              1   2   3   4    5    6   7   8   9   10
rc1    vcc     n01             290
rc2    vcc     n02             290
rc3    vcc     n04             150
q1     n01     in1     n03     2N3904
q2     n01     in2     n03     2N3904
q3     n01     in3     n03     2N3904
q4     n04     n06     n03     2N3904
q5     n04     n06     n05     2N3904
q6     n02     in4     n05     2N3904
q7     n02     in5     n05     2N3904
q8     n02     in6     n05     2N3904
q9     vcc     n08     n07     2N3904
rb1    vcc     n08             300
rb2    n08     n09             2550
d1     n09     n10             1N4148
d2     n10     vee             1N4148
re1    n03     vee             1240
re2    n05     vee             1240
re3    n06     vee             1240
q10    vcc     n02     nor2    2N3904
q11    vcc     n01     nor1    2N3904
ro1    nor1    vee             2000
ro2    nor2    vee             2000
.ends MC312A

.end
