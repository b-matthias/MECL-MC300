MC304.cir
*
* SPICE netlist for the Motorola MC304 ECL circuit
*
* Bias circuit required for other MECL circuits (aka Vbb)
* this circuit is specified to drive up to 25 logic eolements 
* ref page 2-29
*
* Models
*
.import 2N3904.mod
.import 1N4148.mod
*
* Circuit netlist
*
.subckt MC304 vbb  vee  vcc  tp
*             vbb  vee  vcc  tp
r1     vcc     tp              300
q1     vcc     tp      vbb     2N3904
r3     vbb     vee             2000
r2     tp      01              2550
d1     01      02              1N4148
d2     02      vee             1N4148
.ends MC304

.end
