MC352.cir
*
* SPICE netlist for the Motorola MC352 ECL circuit
*
* R-S Flip-Flop, DC coupled with expandable input, and non-buffered output
* ref page 2-52 see also MC352A
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC352 ehi vee vcc nq q set1 set2 elo res1 res2
*             1   2   3   4  5 6    7    8   9    10
rc1    vcc     n01             300
rc2    vcc     ehi             300
q1     vcc     n01     nq      2N3904
q2     vcc     ehi     q       2N3904
q3     n01     set1    elo     2N3904
q4     n01     set2    elo     2N3904
q5     n01     q       n04     2N3904
q6     ehi     nq      n04     2N3904
q7     ehi     res1    elo     2N3904
q8     ehi     res2    elo     2N3904
re1    nq      vee             2000
re2    n04     elo             105
re3    elo     vee             1135
re4    q       vee             2000
.ends MC352

.end
