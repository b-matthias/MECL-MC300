MC305.cir
*
* SPICE netlist for the Motorola MC305 ECL circuit
*
* 5-input expander
* see also MC302, MC306, MC307 and MC315
* ref page 2-28
*
* Models
*
.import 2N3904.mod
*
* Circuit netlist
*
.subckt MC305 nc nc nc elo ehi in1 in2 in3 in4 in5
*             1  2  3  4   5   6   7   8   9   10
q1     ehi     in1     elo     2N3904
q2     ehi     in2     elo     2N3904
q3     ehi     in3     elo     2N3904
q4     ehi     in4     elo     2N3904
q5     ehi     in5     elo     2N3904
.ends MC305

.end
